// Verilog test fixture created from schematic C:\Users\Name\Documents\CS120A\Lab5\FA4Bit_5BitReg.sch - Mon Nov 04 16:32:02 2019

`timescale 1ns / 1ps

module FA4Bit_5BitReg_FA4Bit_5BitReg_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   FA4Bit_5BitReg UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
