`timescale 1ns / 1ps

module FullAdder_FullAdder_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   FullAdder UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
